`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:50:33 12/06/2020 
// Design Name: 
// Module Name:    Year_sep 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Year_sep(NUMBER, N1000, N100, N10, N1);
	input [6:0] NUMBER;
	output [7:0] N10, N1;
	
	reg [3:0] number10, number1;


endmodule
