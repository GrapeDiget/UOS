`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    04:14:51 11/08/2020 
// Design Name: 
// Module Name:    lab_04 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module lab_04(clk_1k, resetn, seg_com, seg_data);
	input clk_1k, resetn;
	output reg [3:0] seg_com;
	output reg [7:0] seg_data;
	
	reg sign = 1'b1; //0: ���, 1: ����
	reg [3:0] hundreds = 4'd1;  //���� �ڸ� bcd
	reg [3:0] tens = 4'd3;      //���� �ڸ� bcd
	reg [3:0] ones = 4'd7;      //���� �ڸ� bcd
	
	wire [7:0] s_segment;
	assign s_segment = sign ? 8'b00000010 : 8'b00000000;  //��ȣ�� fnd ���ڷ� ��ȯ
	wire [7:0] h_segment;
	fnd_decoder U0 (.bcd(hundreds), .out(h_segment));     //bcd�� fnd ���ڷ� ��ȯ
	wire [7:0] t_segment;
	fnd_decoder U1 (.bcd(tens), .out(t_segment));			//bcd�� fnd ���ڷ� ��ȯ
	wire [7:0] o_segment;
	fnd_decoder U2 (.bcd(ones), .out(o_segment));			//bcd�� fnd ���ڷ� ��ȯ
	
	integer CNT_SCAN;
	
	always @(negedge resetn or posedge clk_1k) begin
		if(~resetn)
			CNT_SCAN = 0;
		else begin
			if(CNT_SCAN >= 3)
				CNT_SCAN = 0;
			else
				CNT_SCAN = CNT_SCAN + 1;
		end
	end
	
	always @(negedge resetn or posedge clk_1k) begin
		if(~resetn) begin
			seg_com = 4'hF;
			seg_data = 8'h00;
		end
		else begin
			case (CNT_SCAN)
				0 : begin
					seg_com = 4'b0111;
					seg_data = s_segment;
				end
				1 : begin
					seg_com = 4'b1011;
					seg_data = h_segment;
				end
				2: begin
					seg_com = 4'b1101;
					seg_data = t_segment;
				end
				3 : begin
					seg_com = 4'b1110;
					seg_data = o_segment;
				end
				default : begin
					seg_com = 4'hF;
					seg_data = 8'h00;
				end
			endcase
		end
	end

endmodule
