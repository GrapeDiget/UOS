`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:07:28 12/01/2020 
// Design Name: 
// Module Name:    Time_mode 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Time_mode(RESET, CLK, TIME_DATA);
	input RESET, CLK;
	output [31:0] TIME_DATA;
	
	


endmodule
